LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ROM_S IS
PORT (a: IN STD_LOGIC_VECTOR(3 downto 0);
	  d: OUT STD_LOGIC_VECTOR (7 downto 0)
	  );
END ROM_S;

ARCHITECTURE MEMMATRIX OF ROM_S IS

SIGNAL y: STD_LOGIC_VECTOR (15 downto 0);

BEGIN

WITH a(3 downto 0) SELECT
y<= "1000000000000000" when "0000",
	"0100000000000000" when "0001",
	"0010000000000000" when "0010",
	"0001000000000000" when "0011",
	"0000100000000000" when "0100",
	"0000010000000000" when "0101",
	"0000001000000000" when "0110",
	"0000000100000000" when "0111",
	"0000000010000000" when "1000",
	"0000000001000000" when "1001",
	"0000000000100000" when "1010",
	"0000000000010000" when "1011",
	"0000000000001000" when "1100",
	"0000000000000100" when "1101",
	"0000000000000010" when "1110",
	"0000000000000001" when "1111",
	"ZZZZZZZZZZZZZZZZ" when OTHERS;
	
	
WITH y(15 downto 0) SELECT
d<=  "11111111" when "0000000000000001",
	 "00000000" when "0000000000000010", 
	 "10010000" when "0000000000000100",  
	 "00000011" when "0000000000001000",
	 "00001111" when "0000000000010000",
	 "11110000" when "0000000000100000",
	 "00000000" when "0000000001000000", 
	 "00000000" when "0000000010000000",
	 "00000001" when "0000000100000000",
	 "00000010" when "0000001000000000",
	 "00000100" when "0000010000000000",
	 "00001000" when "0000100000000000",
	 "00010000" when "0001000000000000",
	 "00100000" when "0010000000000000",
	 "01000000" when "0100000000000000",
	 "10000000" when "1000000000000000",
	 "ZZZZZZZZ" when OTHERS;

END MEMMATRIX;